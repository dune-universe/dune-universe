package SomePkg;

  localparam IMP_DAT_BITS = 2;
  localparam MOD_BITS = 32'h8;
  localparam BIN_BITS = 32'b1;
  localparam OCT_BITS = 32'o5;

  localparam bit BIT_DAT_BITS = 2;
  localparam bit BIT_MOD_BITS = 32'h8;
  localparam bit BIT_BIN_BITS = 32'b1;
  localparam bit BIT_OCT_BITS = 32'o5;

  localparam logic LOG_DAT_BITS = 2;
  localparam logic LOG_MOD_BITS = 32'h8;
  localparam logic LOG_BIN_BITS = 32'b1;
  localparam logic LOG_OCT_BITS = 32'o5;

  localparam reg REG_DAT_BITS = 2;
  localparam reg REG_MOD_BITS = 32'h8;
  localparam reg REG_BIN_BITS = 32'b1;
  localparam reg REG_OCT_BITS = 32'o5;

  localparam byte BYTE_DAT_BITS = 2;
  localparam byte BYTE_MOD_BITS = 32'h8;
  localparam byte BYTE_BIN_BITS = 32'b1;
  localparam byte BYTE_OCT_BITS = 32'o5;

  localparam shortint SHORTINT_DAT_BITS = 2;
  localparam shortint SHORTINT_MOD_BITS = 32'h8;
  localparam shortint SHORTINT_BIN_BITS = 32'b1;
  localparam shortint SHORTINT_OCT_BITS = 32'o5;

  localparam int INT_DAT_BITS = 2;
  localparam int INT_MOD_BITS = 32'h8;
  localparam int INT_BIN_BITS = 32'b1;
  localparam int INT_OCT_BITS = 32'o5;

  localparam longint LONGINT_DAT_BITS = 2;
  localparam longint LONGINT_MOD_BITS = 32'h8;
  localparam longint LONGINT_BIN_BITS = 32'b1;
  localparam longint LONGINT_OCT_BITS = 32'o5;

  localparam integer INTEGER_DAT_BITS = 2;
  localparam integer INTEGER_MOD_BITS = 32'h8;
  localparam integer INTEGER_BIN_BITS = 32'b1;
  localparam integer INTEGER_OCT_BITS = 32'o5;

  localparam time TIME_DAT_BITS = 2;
  localparam time TIME_MOD_BITS = 32'h8;
  localparam time TIME_BIN_BITS = 32'b1;
  localparam time TIME_OCT_BITS = 32'o5;

endpackage
